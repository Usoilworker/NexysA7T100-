`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/26/2023 10:45:19 PM
// Design Name: 
// Module Name: bramv2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// Single-Port Block RAM Write-First Mode (recommended template)
// File: rams_sp_wf.v
module rams_sp_wf (clk, we, en, addr, di, dout);
input clk;
input we;
input en;
input [15:0] addr;
input [15:0] di;
output [15:0] dout;
reg [15:0] RAM [65535:0];
reg [15:0] dout;

always @(posedge clk)
    begin
        if (en)
        begin
            if (we)
                begin
                RAM[addr] <= di;
                end
             end
            dout <= RAM[addr];
end
endmodule

